module cpu(clk,rst_n,hlt,pc);

input clk;
input rst_n; 
output hlt;
output [15:0] pc;

//todo



endmodule
