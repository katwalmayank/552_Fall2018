module RED_16bit(A, B, Sum);

input [15:0] A, B;
output [15:0] Sum;


endmodule