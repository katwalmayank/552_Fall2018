module RegisterFile(clk,rst,SrcReg1,SrcReg2,DstReg,WriteReg,DstData,SrcData1,SrcData2);

input clk;
input rst;
input [3:0] SrcReg1,SrcReg2; 
input [3:0] DstReg;
input WriteReg;
input [15:0] DstData;
inout [15:0] SrcData1, SrcData2;

//TODO


endmodule

